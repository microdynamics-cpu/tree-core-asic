module S011HD1P_X32Y2D128_BW (
    output reg [     Bits-1:0] Q,
    input                      CLK,
    input                      CEN,
    input                      WEN,
    input      [Wen_Width-1:0] BWEN,
    input      [Add_Width-1:0] A,
    input      [     Bits-1:0] D
);
  localparam Bits = 128;
  localparam Word_Depth = 64;
  localparam Add_Width = 6;
  localparam Wen_Width = 128;

  wire cen = ~CEN;
  wire wen = ~WEN;
  wire [Wen_Width-1:0] bwen = ~BWEN;
  reg  [     Bits-1:0] ram[0:Word_Depth-1];

  always @(posedge CLK) begin
    if (cen && wen) begin
      ram[A] <= (D & bwen) | (ram[A] & ~bwen);
    end
    Q <= cen && !wen ? ram[A] : {4{$random}};
  end

endmodule

module pll
(
    input clk,
    input [2:0] cfg,
    output pll_clk
);

assign pll_clk = clk;

endmodule